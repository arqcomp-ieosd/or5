-- que se terminel anio
